module stalls_hazard(ResultSrcE,RS1_D,RS2_D,RD_E,StallF,StallD,FlushE);

    //Declare I/Os
    input ResultSrcE;
    input [4:0] RD_E;
    input [4:0] RS1_D,RS2_D;
    output StallF,StallD,FlushE;

    //Extract RS1D & RS2D from InstrD
   // wire [4:0] RS1_D = InstrD[19:15];
    //wire [4:0] RS2_D = InstrD[24:20];

    // Compute lwStall based on load word dependency
    wire lwStall;
    //Logic
    assign lwStall = ResultSrcE & ((RS1_D == RD_E) | (RS2_D == RD_E));
    assign StallF = lwStall;
    assign StallD = lwStall;
    assign FlushE = lwStall;
  
endmodule